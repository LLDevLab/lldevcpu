library ieee;
use ieee.std_logic_1164.all;

use work.lldevcpu_pack.all;

entity i2c_master is
	-- data_out - outgoing data
	-- data_in - incoming data 
	port(clk: in std_logic; start: in boolean; addr: in data8; data_out: in data8; sda: inout std_logic := '1'; data_in: out data8 := X"00"; 
			scl: buffer std_logic := '1'; ready: out boolean := true);
end entity;

architecture i2c_master_arch of i2c_master is	
	type bool_arr_2 is array(0 to 1) of boolean;
	
	signal sda_rw_s: i2c_rw := i2c_write;
	signal sda_s: std_logic := '1';
	signal i2c_state_s: i2c_state;
	signal i2c_state_addr_s: i2c_send_state;
	signal i2c_state_data_s: i2c_send_state;
	signal addr_ack_s: std_logic := '1';
	signal data_ack_s: std_logic := '1';
	signal addr_s: data8 := X"00";
	signal data_s: data8 := X"00";
	
	signal sda_ready_s: boolean := true;
	signal scl_ready_s: boolean := true;
	
	function generate_scl(scl_in: std_logic) return std_logic is
	begin
		if(scl_in = '1') then
			return '0';
		else
			return '1';
		end if;
	end generate_scl;
begin
	sda <= sda_s when sda_rw_s = i2c_write else 'Z';
	ready <= sda_ready_s and scl_ready_s;
	
	-- process, that manages i2c states
	state_proc: process(clk, start)
	begin
		if(falling_edge(clk)) then
			case i2c_state_s is
				when i2c_idle =>
					if(start) then
						i2c_state_s <= i2c_start;
						scl_ready_s <= false;
						scl <= '1';
					end if;
				when i2c_start =>
					if(sda = '0' and scl = '0') then
						i2c_state_s <= i2c_addr_send;
						sda_rw_s <= i2c_write;
					elsif(sda = '0' and scl = '1') then
						scl <= '0';
					end if;
				when i2c_addr_send =>
					if(scl = '1') then
						case i2c_state_addr_s is
							when i2c_sending_ack =>
								sda_rw_s <= i2c_read;
							when i2c_sending_rdy =>
								i2c_state_s <= i2c_data_send;
								
								if(addr_s(i2c_addr_rw_bit) = '0') then
									sda_rw_s <= i2c_write;
								else
									sda_rw_s <= i2c_read;
								end if;
							when others =>
								null;
						end case;
					end if;
					
					scl <= generate_scl(scl);
				when i2c_data_send =>
					if(scl = '1') then
						if(addr_s(i2c_addr_rw_bit) = '0') then
							case i2c_state_data_s is
								when i2c_sending =>
									sda_rw_s <= i2c_write;
								when i2c_sending_ack =>
									sda_rw_s <= i2c_read;
								when i2c_sending_rdy =>
									i2c_state_s <= i2c_stop;
									sda_rw_s <= i2c_write;
								when others =>
									null;
							end case;
						else
							case i2c_state_data_s is
								when i2c_sending =>
									sda_rw_s <= i2c_read;
								when i2c_sending_ack =>
									sda_rw_s <= i2c_write;
								when i2c_sending_rdy =>
									i2c_state_s <= i2c_stop;
									sda_rw_s <= i2c_write;
								when others =>
									null;
							end case;
						end if;
					end if;

					scl <= generate_scl(scl);
				when i2c_stop =>
					scl <= '1';
					if(sda_s = '1') then
						i2c_state_s <= i2c_idle;
						scl_ready_s <= true;
					end if;
				when others =>
					null;
			end case;
		end if;
	end process state_proc;
	
	sda_proc: process(clk)
		variable cnt_v: data8_range := 0;
	begin
		if(rising_edge(clk)) then
			case i2c_state_s is
				when i2c_start =>
					data_s <= data_out;
					addr_s <= addr;
					sda_s <= '0';
					sda_ready_s <= false;
					i2c_state_addr_s <= i2c_sending;
					i2c_state_data_s <= i2c_sending;
				when i2c_addr_send =>
					case i2c_state_addr_s is
						when i2c_sending =>
							if(scl = '0') then
								sda_s <= addr_s(cnt_v);
							else
								if(cnt_v < 7) then
									cnt_v := cnt_v + 1;
								else
									cnt_v := 0;
									i2c_state_addr_s <= i2c_sending_ack;
								end if;
							end if;
						when i2c_sending_ack =>
							if(scl = '1') then
								addr_ack_s <= sda;
								i2c_state_addr_s <= i2c_sending_rdy;
							end if;
						when others =>
							null;
					end case;
				when i2c_data_send =>
					if(addr_s(i2c_addr_rw_bit) = '0') then
						case i2c_state_data_s is
							when i2c_sending =>
								if(scl = '0') then
									sda_s <= data_s(cnt_v);
								else
									if(cnt_v < 7) then
										cnt_v := cnt_v + 1;
									else
										cnt_v := 0;
										i2c_state_data_s <= i2c_sending_ack;
									end if;
								end if;
							when i2c_sending_ack =>
								if(scl = '1') then
									sda_s <= '0';											-- reset sda_s, just in case
									data_ack_s <= sda;
									
									i2c_state_data_s <= i2c_sending_rdy;
								end if;
							when others =>
								null;
						end case;
					else
						case i2c_state_data_s is
							when i2c_sending =>
								if(scl = '1') then
									sda_s <= '0';											-- reset sda_s, just in case
									data_s(cnt_v) <= sda;
									
									if(cnt_v < 7) then
										cnt_v := cnt_v + 1;
									else
										cnt_v := 0;
										i2c_state_data_s <= i2c_sending_ack;
									end if;
								end if;
							when i2c_sending_ack =>
								if(scl = '0') then
									sda_s <= '0';
								else
									i2c_state_data_s <= i2c_sending_rdy;
								end if;
							when others =>
								null;
						end case;
					end if;
				when i2c_stop =>
					if(scl = '1') then
						sda_s <= '1';
					end if;
					
					data_in <= data_s;					
					sda_ready_s <= true;
				when others =>
					null;
			end case;
		end if;
	end process sda_proc;
end i2c_master_arch;